localparam [4:0] ADD_OP = 5'b01001;
localparam [4:0] SUB_OP = 5'b00110;
localparam [4:0] A_PLUS_A_AND_B_OP = 5'b01000;
localparam [4:0] A_PLUS_A_OP = 5'b01100;
localparam [4:0] AND_OP = 5'b11011;
localparam [4:0] OR_OP = 5'b11110;
localparam [4:0] XOR_OP = 5'b10110;
localparam [4:0] INV_B_OP = 5'b10101;